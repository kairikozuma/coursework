// UCDB API User Guide Example
//
// Copyright 2013 Mentor Graphics Corporation
//
// All Rights Reserved.
//
// THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION WHICH IS THE
// PROPERTY OF MENTOR GRAPHICS CORPORATION OR ITS LICENSORS AND IS SUBJECT TO
// LICENSE TERMS.

module top;
    enum { a, b, c } t = a;
    initial begin
        #1; t = c;
        #1; t = b;
    end
endmodule
